-------------------------------------------------------------------------------
--
-- Title       : 
-- Design      : lab_10_11
-- Author      : 
-- Company     : 
--
-------------------------------------------------------------------------------
--
-- File        : C:\Users\Hubert Jarosz\Documents\GitHub\UniwersytetZielonogorski\UkladyCyfrowe\Lab_10-11\Lab_10_11\lab_10_11\compile\Zad_06.vhd
-- Generated   : Mon Jan 20 10:22:47 2025
-- From        : C:\Users\Hubert Jarosz\Documents\GitHub\UniwersytetZielonogorski\UkladyCyfrowe\Lab_10-11\Lab_10_11\lab_10_11\src\Zad_06\Zad_06.bde
-- By          : Bde2Vhdl ver. 2.6
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------
-- Design unit header --
library IEEE;
use IEEE.std_logic_1164.all;

entity Zad_06 is
  port(
       X : in STD_LOGIC;
       Clock : in STD_LOGIC;
       Reset : in STD_LOGIC;
       Y2 : buffer STD_LOGIC;
       Y1 : buffer STD_LOGIC;
       Y0 : buffer STD_LOGIC
  );
end Zad_06;

architecture Zad_06 of Zad_06 is

begin

end Zad_06;
